LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY mux_4a1_M IS
generic ( n: integer:=4);
PORT(DIN:IN STD_LOGIC_VECTOR(n-1 DOWNTO 0);
SEL:IN STD_LOGIC_VECTOR(1 DOWNTO 0);DOUT:OUT STD_LOGIC);
END mux_4a1_M  ;
ARCHITECTURE BEH123 OF mux_4a1_M  IS
BEGIN
PROCESS(DIN,SEL)
BEGIN
CASE SEL IS
WHEN"00"=>DOUT<=DIN(0);
WHEN"01"=>DOUT<=DIN(1);
WHEN"10"=>DOUT<=DIN(2);
WHEN"11"=>DOUT<=DIN(3);
WHEN OTHERS=>DOUT<='Z';
END CASE;
END PROCESS;
END BEH123;