LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY mux_8a1 IS
generic ( n: integer:=8);
PORT(DIN:IN STD_LOGIC_VECTOR(n-1 DOWNTO 0);
SEL:IN STD_LOGIC_VECTOR(2 DOWNTO 0);DOUT:OUT STD_LOGIC);
END mux_8a1 ;
ARCHITECTURE BEH123 OF mux_8a1 IS
BEGIN
PROCESS(DIN,SEL)
BEGIN
CASE SEL IS
WHEN"000"=>DOUT<=DIN(0);
WHEN"001"=>DOUT<=DIN(1);
WHEN"010"=>DOUT<=DIN(2);
WHEN"011"=>DOUT<=DIN(3);
WHEN"100"=>DOUT<=DIN(4);
WHEN"101"=>DOUT<=DIN(5);
WHEN"110"=>DOUT<=DIN(6);
WHEN"111"=>DOUT<=DIN(7);
WHEN OTHERS=>DOUT<='Z';
END CASE;
END PROCESS;
END BEH123;